module main
(
);

//

endmodule
