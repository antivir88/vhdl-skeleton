module vidac
(
);

//

endmodule
